* C:\FOSSEE\eSim\library\SubcircuitLibrary\HA_test\HA_test.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 6/11/2024 6:43:09 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M3  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M3-Pad3_ Net-_M3-Pad3_ eSim_MOS_P		
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ GND GND eSim_MOS_N		
M4  Net-_M2-Pad1_ Net-_M1-Pad2_ GND Net-_M3-Pad3_ eSim_MOS_P		
M2  Net-_M2-Pad1_ Net-_M1-Pad2_ /B GND eSim_MOS_N		
M6  /Sum /B Net-_M1-Pad2_ Net-_M3-Pad3_ eSim_MOS_P		
M5  /Sum /B Net-_M1-Pad1_ GND eSim_MOS_N		
v1  Net-_M3-Pad3_ GND DC		
U1  Net-_M1-Pad2_ /B /Sum Net-_M2-Pad1_ PORT		

.end
