* C:\FOSSEE\eSim\library\SubcircuitLibrary\FA_test\FA_test.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 6/11/2024 8:02:28 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M1  Net-_M1-Pad1_ /A /B /VDD eSim_MOS_P		
M2  Net-_M1-Pad1_ /A Net-_M2-Pad3_ GND eSim_MOS_N		
M6  /C Net-_M1-Pad1_ Net-_M6-Pad3_ GND eSim_MOS_N		
M3  Net-_M2-Pad3_ /B GND GND eSim_MOS_N		
M7  Net-_M6-Pad3_ /C GND GND eSim_MOS_N		
M4  Net-_M1-Pad1_ /B /A /VDD eSim_MOS_P		
M5  /C Net-_M1-Pad1_ /C /VDD eSim_MOS_P		
M8  /C /C Net-_M1-Pad1_ /VDD eSim_MOS_P		
v1  /VDD GND DC		
U1  /A /B /C /C /C PORT		

.end
