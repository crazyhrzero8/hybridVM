* C:\FOSSEE\eSim\library\SubcircuitLibrary\and_test\and_test.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 8/11/2024 10:22:34 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M1  Net-_M1-Pad1_ /A /VDD /VDD eSim_MOS_P		
M4  Net-_M1-Pad1_ /B /VDD /VDD eSim_MOS_P		
M6  /Y Net-_M1-Pad1_ /VDD /VDD eSim_MOS_P		
M2  Net-_M1-Pad1_ /A Net-_M2-Pad3_ GND eSim_MOS_N		
M3  Net-_M2-Pad3_ /B GND GND eSim_MOS_N		
M5  /Y Net-_M1-Pad1_ GND GND eSim_MOS_N		
v1  GND /VDD DC		
U1  /A /B /Y PORT		

.end
